package i2cmb_env_pkg;
    import ncsu_pkg::*;
    import i2c_pkg::*;
    import wb_pkg::*;
    import data_types_pkg::*;
    `include "src/i2cmb_generator.svh"
    `include "src/i2cmb_env_configuration.svh"
    `include "src/i2cmb_scoreboard.svh"
    `include "src/i2cmb_predictor.svh"
    `include "src/i2cmb_coverage.svh"
    `include "src/i2cmb_environment.svh"
    `include "src/i2cmb_test.svh"
    `include "src/i2cmb_test_random.svh"
    `include "src/test_i2cmb_reads.svh"
    `include "src/test_i2cmb_writes.svh"
    `include "src/test_i2cmb_reg_addrs.svh"
    `include "src/test_i2cmb_two_starts.svh"
    `include "src/test_i2cmb_two_stops.svh"
    `include "src/test_i2cmb_write_before_data.svh"
    `include "src/test_i2cmb_reg_inits.svh"

endpackage
