class i2c_agent extends ncsu_object;

endclass