class i2cmb_test extends ncsu_component;
    // i2cmb_generator generator;
    // i2cmb_env_configuration configuration;
    // i2cmb_environment environment;

    // function new(string name = "", ncsu_component #(T) parent = null); 
    //     super.new(name,parent);
    //     configuration = new("configuration");
    //     configuration.sample_coverage();
    //     environment = new("environment",this);
    //     environment.set_configuration(configuration);
    //     environment.build();
    //     generator = new("generator",this);
    //     generator.set_agent(environment.get_p0_agent());
    // endfunction

    // virtual task run();
    //     environment.run();
    //     generator.run();
    // endtask
    
endclass