class i2cmb_predictor;

endclass