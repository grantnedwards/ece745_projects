class i2cmb_generator;

endclass