class wb_transaction;


endclass