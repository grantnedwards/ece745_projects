class i2c_driver;

endclass