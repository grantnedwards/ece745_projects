class i2cmb_env_configuration;

endclass