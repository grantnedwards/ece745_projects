class i2c_configuration;

endclass