class i2c_monitor;

endclass