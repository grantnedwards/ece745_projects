class wb_monitor;

endclass