class i2cmb_coverage;

endclass