class i2cmb_scoreboard;

endclass
