class wb_transaction extends ncsu_transaction;


endclass