class wb_agent;

endclass