class i2c_agent;
    virtual i2c_driver driver;
    virtual i2c_monitor monitor;
    
endclass