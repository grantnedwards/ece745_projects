class wb_configuration;

endclass