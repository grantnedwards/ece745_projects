class i2c_agent;

endclass