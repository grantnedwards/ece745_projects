class i2cmb_test;

endclass