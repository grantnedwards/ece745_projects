class i2c_transaction extends ncsu_transaction;

endclass