class wb_driver;

endclass