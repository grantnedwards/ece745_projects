class wb_agent;
    virtual wb_driver driver;
    virtual wb_monitor monitor;

    
endclass