class i2cmb_environment;

endclass