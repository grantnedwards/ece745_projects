class i2c_driver extends ;

endclass