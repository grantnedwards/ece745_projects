class i2cmb_env_configuration extends ncsu_configuration;
    virtual wb_configuration wishbone;
    virtual i2c_configuration i2c;

    
endclass