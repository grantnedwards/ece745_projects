class i2cmb_environment;
    // wb_agent wishbone_side;
    // i2c_agent i2c_side;

    // i2cmb_predictor predictor;
    // i2cmb_coverage coverage;
    // i2cmb_scoreboard scoreboard;
endclass