class i2cmb_test;
    virtual i2cmb_generator generator;
    virtual i2cmb_env_configuration env_config;
    virtual i2cmb_environment environment;
    
endclass