class i2c_transaction;

endclass